package nvme_trans_lib_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;

  `include "nvme_enum_lib.sv"
  `include "nvme_struct_lib.sv"
  `include "identify_controller_data_struct.sv"
endpackage
