package host_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "nvme_macros.svh"

  `include "base_q.svh"
endpackage
