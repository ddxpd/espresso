/************Admin Command Opcode Enum************/
typedef enum {
  DeleteIOSubmissionQueue = 'h00,
  CreateIOSubmissionQueue = 'h01,
  GetLogPage = 'h02,
  DeleteIOCompletionQueue = 'h04,
  CreateIOCompletionQueue = 'h05,
  Identify = 'h06,
  Abort = 'h08,
  SetFeatures = 'h09,
  GetFeatures = 'h0A,
  AsynchronousEventRequest = 'h0C,
  NamespaceManagement = 'h0D,
  FirmwareCommit = 'h10,
  FirmwareImageDownload = 'h11,
  DeviceSelf_test = 'h14,
  NamespaceAttachment = 'h15,
  KeepAlive = 'h18,
  DirectiveSend = 'h19,
  DirectiveReceive = 'h1A,
  VirtualizationManagement = 'h1C,
  NVMeMISend = 'h1D,
  NVMeMIReceive = 'h1E,
  CapacityManagement = 'h20,
  DiscoveryInformationManagement = 'h21,
  FabricZoningReceive = 'h22,
  Lockdown = 'h24,
  FabricZoningLookup = 'h25,
  ClearExportedNVMResourceConfiguration = 'h28,
  FabricZoningSend = 'h29,
  CreateExportedNVMSubsystem = 'h2A,
  ManageExportedNVMSubsystem = 'h2D,
  ManageExportedNamespace = 'h31,
  ManageExportedPort = 'h35,
  SendDiscoveryLogPage = 'h39,
  TrackSend = 'h3D,
  TrackReceive = 'h3E,
  MigrationSend = 'h41,
  MigrationReceive = 'h42,
  ControllerDataQueue = 'h45,
  DoorbellBufferConfig = 'h7C,
  FabricsCommands = 'h7F,
  FormatNVM = 'h80,
  SecuritySend = 'h81,
  SecurityReceive = 'h82,
  Sanitize = 'h84,
  LoadProgram = 'h85,
  GetLBAStatus = 'h86,
  ProgramActivationManagement = 'h88,
  MemoryRangeSetManagement = 'h89
  //Vendorspecific = 'hC0h to FF,
} E_ADMIN_CMD_OPCODE;


/*****************GET FEATURE  FEATURE ID********************/
typedef enum {
  Arbitration = 'h01, 
  PowerManagement = 'h02, 
  TemperatureThreshold = 'h04, 
  VolatileWriteCache = 'h06, 
  NumberofQueues = 'h07, 
  InterruptCoalescing = 'h08, 
  InterruptVectorConfiguration = 'h09, 
  AsynchronousEventConfiguration = 'h0B, 
  AutonomousPowerStateTransition = 'h0C, 
  HostMemoryBuffer = 'h0D, 
  Timestamp = 'h0E, 
  KeepAliveTimer = 'h0F, 
  HostControlledThermalManagement = 'h10, 
  NonOperationalPowerStateConfig = 'h11, 
  ReadRecoveryLevelConfig = 'h12, 
  PredictableLatencyModeConfig = 'h13, 
  PredictableLatencyModeWindow = 'h14, 
  HostBehaviorSupport = 'h16, 
  SanitizeConfig = 'h17, 
  EnduranceGroupEventConfiguration = 'h18, 
  IOCommandSetProfile = 'h19, 
  SpinupControl = 'h1A, 
  PowerLossSignalingConfig = 'h1B, 
  FlexibleDataPlacement = 'h1D, 
  FlexibleDataPlacementEvents = 'h1E, 
  NamespaceAdminLabel = 'h1F, 
  ControllerDataQueueID = 'h21, 
  EmbeddedManagementControllerAddress = 'h78, 
  HostManagementAgentAddress = 'h79, 
  EnhancedControllerMetadata = 'h7D, 
  ControllerMetadata = 'h7E, 
  NamespaceMetadata = 'h7F, 
  SoftwareProgressMarker = 'h80, 
  HostIdentifier = 'h81, 
  ReservationNotificationMask = 'h82, 
  ReservationPersistence = 'h83, 
  NamespaceWriteProtectionConfig = 'h84, 
  BootPartitionWriteProtectionConfig = 'h85 
} E_GET_FEATURE_FEATURE_ID;


/*****************GET LOG PAGE  PAGE ID********************/
typedef enum {
  SupportedLogPages = 'h00, 
  ErrorInformation = 'h01, 
  ControllerNamespace = 'h02, 
  FirmwareSlotInformation = 'h03, 
  ChangedAttachedNamespaceList = 'h04, 
  CommandsSupportedandEffects = 'h05, 
  DeviceSelftest = 'h06, 
  TelemetryHost_Initiated = 'h07, 
  TelemetryControllerInitiated = 'h08, 
  EnduranceGroupInformation = 'h09, 
  PredictableLatencyPerNVMSet = 'h0A, 
  PredictableLatencyEventAggregate = 'h0B, 
  AsymmetricNamespaceAccess = 'h0C, 
  PersistentEventLog = 'h0D, 
  EnduranceGroupEventAggregate = 'h0F, 
  DomainNVMsubsystem = 'h10, 
  SupportedCapacityConfigurationList = 'h11, 
  FeatureIdentifiersSupportedandEffects = 'h12, 
  NVMeMICommandsSupportedandEffects = 'h13, 
  CommandandFeatureLockdown = 'h14, 
  BootPartition = 'h15, 
  RotationalMediaInformation = 'h16, 
  DispersedNamespaceParticipatingNVMSubsystems = 'h17, 
  ManagementAddressList = 'h18, 
  ReachabilityGroups = 'h1A, 
  ReachabilityAssociations = 'h1B, 
  ChangedAllocatedNamespaceList = 'h1C, 
  FDPConfigurations = 'h20, 
  ReclaimUnitHandleUsage = 'h21, 
  FDPStatistics = 'h22, 
  FDPEvents = 'h23, 
  Discovery = 'h70, 
  HostDiscovery = 'h71, 
  AVEDiscovery = 'h72, 
  PullModelDDCRequest = 'h73, 
  ReservationNotification = 'h80, 
  SanitizeStatus = 'h81 
} E_LOG_PAGE_ID;

typedef enum {
  IdentifyNamespacedatastructure = 'h00, 
  IdentifyControllerdatastructure = 'h01, 
  ActiveNamespaceIDlist = 'h02, 
  NamespaceIdentificationDescriptorlist = 'h03, 
  AnNVMSetList = 'h04, 
  IOCommandSetspecificIdentifyNamespacedatastructure = 'h05, 
  IOCommandSetspecificIdentifyControllerdatastructure = 'h06, 
  ActiveNamespaceIDlistwithIOCommandSet = 'h07, 
  IOCommandSetIndependentIdentifyNamespacedatastructure = 'h08, 
  IdentifyNamespacedatastructureforFormatIndex = 'h09, 
  IOCommandSetspecificIdentifyNamespacedatastructureforFormatIndex = 'h0A, 
  AllocatedNamespaceIDlist = 'h10, 
  IdentifyNamespacedatastructureforallocatedNSID = 'h11, 
  ControllerListofcontrollersattachedtothespecifiedNSID = 'h12, 
  ControllerListofcontrollersthatexistintheNVMsubsystem = 'h13, 
  PrimaryControllerCapabilitiesdatastructure = 'h14, 
  SecondaryControllerlistofcontroller = 'h15, 
  ANamespaceGranularityList = 'h16, 
  AUUIDList = 'h17, 
  DomainList = 'h18, 
  EnduranceGroupList = 'h19, 
  IOCommandSetspecificAllocatedNamespaceIDlist = 'h1A, 
  IOCommandSetspecificIdentifyNamespacedatastructureforAllocatedID = 'h1B, 
  IOCommandSetdatastructure = 'h1C, 
  GetUnderlyingNamespaceList = 'h1D, 
  GetPortsList = 'h1E, 
  IOCommandSetIndependentIdentifyNamespacedatastructureforallocatedNSID = 'h1F, 
  SupportedControllerStateFormats = 'h20 
} E_IDENTIFY_CNS;

typedef enum {
  NVMCommandSet = 'h00, 
  KeyValueCommandSet = 'h01, 
  ZonedNamespaceCommandSet = 'h02, 
  SubsystemLocalMemoryCommandSet = 'h03, 
  ComputationalProgramsCommandSet = 'h04
} E_IDENTIFY_CMD_SET_ID;

/************Completion Status Code Enum************/
typedef enum {
  GenericCommandStatus = 'h0,
  CommandSpecificStatus = 'h1,
  MediaandDataIntegrityErrors = 'h2,
  PathRelatedStatus = 'h3,
  VendorSpecific = 'h7
} E_STATUS_CODE_TYPE;

typedef enum {
  SuccessfulCompletion = 'h00,
  InvalidCommandOpcode = 'h01,
  InvalidFieldinCommand = 'h02,
  CommandIDConflict = 'h03,
  DataTransferError = 'h04,
  CommandsAbortedduetoPowerLossNotification = 'h05,
  InternalError = 'h06,
  CommandAbortRequested = 'h07,
  CommandAbortedduetoSQDeletion = 'h08,
  CommandAbortedduetoFailedFusedCommand = 'h09,
  CommandAbortedduetoMissingFusedCommand = 'h0A,
  InvalidNamespaceorFormat = 'h0B,
  CommandSequenceError = 'h0C,
  InvalidSGLSegmentDescriptor = 'h0D,
  InvalidNumberofSGLDescriptors = 'h0E,
  DataSGLLengthInvalid = 'h0F,
  MetadataSGLLengthInvalid = 'h10,
  SGLDescriptorTypeInvalid = 'h11,
  InvalidUseofControllerMemoryBuffer = 'h12,
  PRPOffsetInvalid = 'h13,
  AtomicWriteUnitExceeded = 'h14,
  OperationDenied = 'h15,
  SGLOffsetInvalid = 'h16,
  Reserved = 'h17,
  HostIdentifierInconsistentFormat = 'h18,
  KeepAliveTimerExpired = 'h19,
  KeepAliveTimeoutInvalid = 'h1A,
  CommandAbortedduetoPreemptandAbort = 'h1B,
  SanitizeFailed = 'h1C,
  SanitizeInProgress = 'h1D,
  SGLDataBlockGranularityInvalid = 'h1E,
  CommandNotSupportedforQueueinCMB = 'h1F,
  NamespaceisWriteProtected = 'h20,
  CommandInterrupted = 'h21,
  TransientTransportError = 'h22,
  CommandProhibitedbyCommandandFeatureLockdown = 'h23,
  AdminCommandMediaNotReady = 'h24,
  InvalidKeyTag = 'h25,
  HostDispersedNamespaceSupportNotEnabled = 'h26,
  HostIdentifierNotInitialized = 'h27,
  IncorrectKey = 'h28,
  FDPDisabled = 'h29,
  InvalidPlacementHandleList = 'h2A,
  LBAOutofRange = 'h80,
  CapacityExceeded = 'h81,
  NamespaceNotReady = 'h82,
  ReservationConflict = 'h83,
  FormatInProgress = 'h84,
  InvalidValueSize = 'h85,
  InvalidKeySize = 'h86,
  KVKeyDoesNotExist = 'h87,
  UnrecoveredError = 'h88,
  KeyExists = 'h89
  //90h to BF, Reserved
  //C0h to FF, Vendor Specific
} E_GENERIC_STATUS_CODE;


typedef enum {
  CompletionQueueInvalid = 'h00,
  InvalidQueueIdentifier = 'h01,
  InvalidQueueSize = 'h02,
  AbortCommandLimitExceeded = 'h03,
  AsynchronousEventRequestLimitExceeded = 'h05,
  InvalidFirmwareSlot = 'h06,
  InvalidFirmwareImage = 'h07,
  InvalidInterruptVector = 'h08,
  InvalidLogPage = 'h09,
  InvalidFormat = 'h0A,
  FirmwareActivationRequiresConventionalReset = 'h0B,
  InvalidQueueDeletion = 'h0C,
  FeatureIdentifierNotSaveable = 'h0D,
  FeatureNotChangeable = 'h0E,
  FeatureNotNamespaceSpecific = 'h0F,
  FirmwareActivationRequiresNVMSubsystemReset = 'h10,
  FirmwareActivationRequiresControllerLevelReset = 'h11,
  FirmwareActivationRequiresMaximumTimeViolation = 'h12,
  FirmwareActivationProhibited = 'h13,
  OverlappingRange = 'h14,
  NamespaceInsufficientCapacity = 'h15,
  NamespaceIdentifierUnavailable = 'h16,
  NamespaceAlreadyAttached = 'h18,
  NamespaceIsPrivate = 'h19,
  NamespaceNotAttached = 'h1A,
  ThinProvisioningNotSupported = 'h1B,
  ControllerListInvalid = 'h1C,
  DeviceSelftestInProgress = 'h1D,
  BootPartitionWriteProhibited = 'h1E,
  InvalidControllerIdentifier = 'h1F,
  InvalidSecondaryControllerState = 'h20,
  InvalidNumberofControllerResources = 'h21,
  InvalidResourceIdentifier = 'h22,
  SanitizeProhibitedWhilePersistentMemoryRegionisEnabled = 'h23,
  ANAGroupIdentifierInvalid = 'h24,
  ANAAttachFailed = 'h25,
  InsufficientCapacity = 'h26,
  NamespaceAttachmentLimitExceeded = 'h27,
  ProhibitionofCommandExecutionNotSupported = 'h28,
  IOCommandSetNotSupported = 'h29,
  IOCommandSetNotEnabled = 'h2A,
  IOCommandSetCombinationRejected = 'h2B,
  InvalidIOCommandSet = 'h2C,
  IdentifierUnavailable = 'h2D,
  NamespaceIsDispersed = 'h2E,
  InvalidDiscoveryInformation = 'h2F,
  ZoningDataStructureLocked = 'h30,
  ZoningDataStructureNotFound = 'h31,
  InsufficientDiscoveryResources = 'h32,
  RequestedFunctionDisabled = 'h33,
  ZoneGroupOriginatorInvalid = 'h34,
  InvalidHost = 'h35,
  InvalidNVMSubsystem = 'h36,
  InvalidControllerDataQueue = 'h37,
  NotEnoughResources = 'h38,
  ControllerSuspended = 'h39,
  ControllerNotSuspended = 'h3A,
  ControllerDataQueueFull = 'h3B
} E_COMMAND_SPECIFIC_STATUS_CODE;


typedef enum {
  CAP_CAP       = 0,
  CAP_VERSION   = 2,
  CAP_INTMS     = 3,
  CAP_INTMC     = 4,
  CAP_CC        = 5,
  CAP_CSTS      = 7,
  CAP_NSSR      = 8,
  CAP_AQA       = 9,
  CAP_ASQ       = 10,
  CAP_ACQ       = 12,
  CAP_CMBLOC    = 14,
  CAP_CMBSZ     = 15,
  CAP_BPINFO    = 16,
  CAP_BPRSEL    = 17,
  CAP_BPMBL     = 18,
  CAP_CMBMSC    = 20,
  CAP_CMBSTS    = 22,
  CAP_CMBEBS    = 23,
  CAP_CMBSWTP   = 24,
  CAP_NSSD      = 25,
  CAP_CRTO      = 26,
  CAP_PMRCAP    = 896,
  CAP_PMRCTL    = 897,
  CAP_PMRSTS    = 898,
  CAP_PMREBS    = 899,
  CAP_PMRSWTP   = 900,
  CAP_PMRMSCL   = 901,
  CAP_PMRMSCU   = 902
} E_CAP_POS;

