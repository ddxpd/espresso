package bfm_pkg;
  import misc_pkg::*;
  `include "host_if.svh"
endpackage
