package misc_pkg;
  `include "nvme_macros.svh"
endpackage
