package host_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;
  import bfm_pkg::*;
  import host_mem_pkg::*;

  `include "base_q.svh"
  `include "nvme_mgr.svh"
  `include "nvme_cmd.svh"
  `include "nvme_cpl_entry.svh"
  `include "dut.svh"
  `include "esp_host_software.svh"
  
  
endpackage

