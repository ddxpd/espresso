package misc_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "nvme_macros.svh"
  `include "nvme_misc.svh"

endpackage
