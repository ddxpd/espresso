package test_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;
  import bfm_pkg::*;
  import host_pkg::*;
  import host_mem_pkg::*;
  import nvme_trans_lib_pkg::*;

  `include "init_test.sv"
  `include "base_test.svh"
  `include "demo_test.sv"
endpackage
