package misc_pkg;
  `include "nvme_macros.svh"
  `include "nvme_misc.svh"

endpackage
