parameter  NUM_DW_SQE = 16;
parameter  NUM_DW_CDE = 4;
parameter  HOST_AXI_WIDTH = 64;


typedef bit[63:0]  U64;
typedef bit[31:0]  U32;
typedef bit[15:0]  U16;
typedef bit[ 7:0]  U8;
