package host_mem_pkg;
  import misc_pkg::*;

  `include "host_memory.svh"
endpackage
