package host_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  
  `include "nvme_macros.svh"

  import test_pkg::*;

  `include "base_q.svh"
  `include "esp_host_software.svh"
  `include "nvme_cmd.svh"
  `include "dut.svh"
  `include "nvme_cpl_entry.svh"
  `include "nvme_mgr.svh"
endpackage

