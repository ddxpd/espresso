package test_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import host_pkg::*;
  `include "init_test.sv"
endpackage
