package host_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;
  import bfm_pkg::*;

  `include "nvme_cmd.svh"
  `include "nvme_cpl_entry.svh"
  `include "nvme_mgr.svh"
  `include "base_q.svh"
  `include "esp_host_software.svh"
  `include "dut.svh"
  
endpackage

