package bfm_pkg;
  import misc_pkg::*;
  typedef virtual host_intf host_vif;
endpackage
