package test_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;
  import bfm_pkg::*;
  import host_pkg::*;
  import host_mem_pkg::*;

  `include "init_test.sv"
  `include "base_test.svh"
endpackage
