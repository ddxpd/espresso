package host_mem_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import misc_pkg::*;

  `include "host_memory.svh"
  `include "host_memory_manager.svh"
endpackage
